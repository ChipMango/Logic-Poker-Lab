
//------------------------------------------------------------------------------
// File Name: test_player_interface.sv
// Description:  Testbench for simulating the player interface and verifying the handshake and command transactions.
// Author: <Student Name>
// Date: <Date>
// Version: 1.0
// Project: ChipMango Lab 03 - Digitally Representing Poker Cards
// License: ChipMango Confidential - For educational purposes only
//------------------------------------------------------------------------------
// Revision History:
//   v1.0 - 07/06/25: Initial file created with module template
//------------------------------------------------------------------------------
