
//------------------------------------------------------------------------------
// File Name:player_fsm_controller.sv
// Description:player interface module that integrates memory, evaluator, and command generator with the FSM.
// Author: <Student Name>
// Date: <Date>
// Version: 1.0
// Project: ChipMango Lab 04 - Digitally Representing Poker Cards
// License: ChipMango Confidential - For educational purposes only
//------------------------------------------------------------------------------
// Revision History:
//   v1.0 - 07/06/25: Initial file created with module template
//------------------------------------------------------------------------------
