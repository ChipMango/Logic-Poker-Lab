
//------------------------------------------------------------------------------
// File Name: test_full_player.sv
// Description:   Testbench for simulating the full player behavior.
// Author: <Student Name>
// Date: <Date>
// Version: 1.0
// Project: ChipMango Lab 06 - Digitally Representing Poker Cards
// License: ChipMango Confidential - For educational purposes only
//------------------------------------------------------------------------------
// Revision History:
//   v1.0 - 08/06/25: Initial file created with module template
//------------------------------------------------------------------------------
