//------------------------------------------------------------------------------
// File Name: test_hand_rank_evaluator.sv
// Description:  Testbench that applies various test cases to the hand evaluator.
// Author: <Student Name>
// Date: <Date>
// Version: 1.0
// Project: ChipMango Lab 01 - Digitally Representing Poker Cards
// License: ChipMango Confidential - For educational purposes only
//------------------------------------------------------------------------------
// Revision History:
//   v1.0 - 06/06/25: Initial file created with module template
//------------------------------------------------------------------------------
