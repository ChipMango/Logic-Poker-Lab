//------------------------------------------------------------------------------
// File Name: personality_lfsr.sv
// Description: Verilog file that implements the LFSR logic to select personalities.
// Author: <Student Name>
// Date: <Date>
// Version: 1.0
// Project: ChipMango Lab 05 - Digitally Representing Poker Cards
// License: ChipMango Confidential - For educational purposes only
//------------------------------------------------------------------------------
// Revision History:
//   v1.0 - 07/06/25: Initial file created with module template
//------------------------------------------------------------------------------
