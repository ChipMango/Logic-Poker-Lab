
//------------------------------------------------------------------------------
// File Name: command_generator.sv
// Description:   module that implements the handshke and command generation.
// Author: <Student Name>
// Date: <Date>
// Version: 1.0
// Project: ChipMango Lab 03 - Digitally Representing Poker Cards
// License: ChipMango Confidential - For educational purposes only
//------------------------------------------------------------------------------
// Revision History:
//   v1.0 - 07/06/25: Initial file created with module template
//------------------------------------------------------------------------------

module command_generator (
 // input  logic        clk,
 // input  logic        rst_n,
 // input  logic [2:0]  action_code, // command to send
//  input  logic        trigger,     // pulse to initiate command
//  output logic [2:0]  cr_cmd,
 // output logic        cr_cmdvld,
//  input  logic        cr_ack,
//  output logic        cmd_done     // pulses when ack received
);

//module body (declarations, logic)


// ...other logic, submodule instantiation



endmodule  // command genearator 









