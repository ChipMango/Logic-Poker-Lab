//------------------------------------------------------------------------------
// File Name: test_game_fsm.sv
// Description: Testbench for simulating the FSM and verifying the state transitions and game flow.
// Author: <Student Name>
// Date: <Date>
// Version: 1.0
// Project: ChipMango Lab 04 - Digitally Representing Poker Cards
// License: ChipMango Confidential - For educational purposes only
//------------------------------------------------------------------------------
// Revision History:
//   v1.0 - 07/06/25: Initial file created with module template
//------------------------------------------------------------------------------

